-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Tue Oct 22 17:06:24 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY control_motor IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clk : IN STD_LOGIC;
        Muro : IN STD_LOGIC := '0';
        MD : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
        MI : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
    );
END control_motor;

ARCHITECTURE BEHAVIOR OF control_motor IS
    TYPE type_fstate IS (Derecho_giroDer,Gira_Der_90,Gira_Izq_90,Derecho_giroIzq);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clk,reg_fstate)
    BEGIN
        IF (clk='1' AND clk'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,Muro)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Derecho_giroDer;
            MD <= "00";
            MI <= "00";
        ELSE
            MD <= "00";
            MI <= "00";
            CASE fstate IS
                WHEN Derecho_giroDer =>
                    IF ((Muro = '1')) THEN
                        reg_fstate <= Gira_Izq_90;
                    ELSIF ((Muro = '0')) THEN
                        reg_fstate <= Derecho_giroDer;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Derecho_giroDer;
                    END IF;

                    MI <= "01";

                    MD <= "01";
                WHEN Gira_Der_90 =>
                    IF ((Muro = '0')) THEN
                        reg_fstate <= Derecho_giroDer;
                    ELSIF ((Muro = '1')) THEN
                        reg_fstate <= Gira_Der_90;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Gira_Der_90;
                    END IF;

                    MI <= "01";

                    MD <= "10";
                WHEN Gira_Izq_90 =>
                    IF ((Muro = '1')) THEN
                        reg_fstate <= Gira_Izq_90;
                    ELSIF ((Muro = '0')) THEN
                        reg_fstate <= Derecho_giroIzq;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Gira_Izq_90;
                    END IF;

                    MI <= "10";

                    MD <= "01";
                WHEN Derecho_giroIzq =>
                    IF ((Muro = '1')) THEN
                        reg_fstate <= Gira_Der_90;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Derecho_giroIzq;
                    END IF;

                    MI <= "01";

                    MD <= "01";
                WHEN OTHERS => 
                    MD <= "XX";
                    MI <= "XX";
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
