library verilog;
use verilog.vl_types.all;
entity Prueba_giros_vlg_vec_tst is
end Prueba_giros_vlg_vec_tst;
